package data_types is
    type array_of_integers is array(integer range <>) of integer;
end package;

